-- Copyright (c) 2025 Chair for Chip Design for Embedded Computing,
--                    TU Braunschweig, Germany
--                    www.tu-braunschweig.de/en/eis
--
-- Use of this source code is governed by an MIT-style
-- license that can be found in the LICENSE file or at
-- https://opensource.org/licenses/MIT.


library ieee;
use ieee.std_logic_1164.all;

use work.aux_pkg.all;

entity nano_imem is
  generic(DEPTH      : natural;
          DEPTH_LOG2 : natural;
          WIDTH_BITS : natural
         );
  port(clk1_i  : in  std_logic;
       clk2_i  : in  std_logic;
       oe_i    : in  std_logic;
       we_i    : in  std_logic;
       addr_i  : in  std_logic_vector(DEPTH_LOG2-1 downto 0);
       -- !! changed for MEH ASIC flashloader with 8 bit load, load 2 4-bit instructions parallel !!
       instr_i : in  std_logic_vector(2*WIDTH_BITS-1 downto 0);  --(WIDTH_BITS-1 downto 0);
       -- !! change end !!
       instr_o : out std_logic_vector(WIDTH_BITS-1 downto 0)
      );
end entity nano_imem;

-- pragma translate_off
use work.nano_rom_image.all; -- this file is generated by the assembler

library top_level;

architecture sync_rom of nano_imem is
  
  component clkgate is
    port(clk : in  std_logic;
         en  : in  std_logic;
         gck : out std_logic);
  end component;
  
  -- MEM Array
  type imem_t is array (0 to DEPTH-1) of std_logic_vector(WIDTH_BITS-1 downto 0);
  
  -- Init Function
  function init_imem(init : image_t) return imem_t is
    variable mem_v : imem_t;
  begin
    for i in 0 to DEPTH-1 loop
        mem_v(i) := init(i)(WIDTH_BITS-1 downto 0);
    end loop; -- i
    return mem_v;
  end function init_imem;
  
  -- ROM Image
  constant imem : imem_t := init_imem(init_image);
  
  -- Address Latch Signals
  signal addr : std_logic_vector(DEPTH_LOG2-1 downto 0);
  
  -- Clock Gating Signals
  signal clk1_oe_gated : std_logic;
  
begin
  
  -- Clock Gating (global output enable)
  clk1_oe_gate : clkgate
    port map(clk => clk1_i,
             en  => oe_i,
             gck => clk1_oe_gated);
  
  -- Address Latch
  addr_lat : process(oe_i, addr_i)
  begin
    if oe_i = '1' then
      addr <= addr_i;
    end if;
  end process addr_lat;
  
  -- Output Mux
  out_mux : process(clk1_oe_gated)
    variable dvec : std_logic_vector((2**DEPTH_LOG2)*WIDTH_BITS-1 downto 0);
    variable dout : std_logic_vector(WIDTH_BITS-1                 downto 0);
  begin
    if rising_edge(clk1_oe_gated) then
      dvec := (others => '-');
      for i in 0 to DEPTH-1 loop
        dvec((i+1)*WIDTH_BITS-1 downto i*WIDTH_BITS) := imem(i);
      end loop; --i
      dout := muxtree(dvec, addr, WIDTH_BITS);
      instr_o <= dout;
    end if;
  end process out_mux;
  
end architecture sync_rom;
-- pragma translate_on
