-- Copyright (c) 2022 Chair for Chip Design for Embedded Computing,
--                    Technische Universitaet Braunschweig, Germany
--                    www.tu-braunschweig.de/en/eis
--
-- Use of this source code is governed by an MIT-style
-- license that can be found in the LICENSE file or at
-- https://opensource.org/licenses/MIT.


package func_pkg is

  -- RTC
  constant FUNC_RTC_CNT_W_C : natural := 17;  -- Width of RTC counter
  
end package func_pkg;
