-- Copyright (c) 2025 Chair for Chip Design for Embedded Computing,
--                    TU Braunschweig, Germany
--                    www.tu-braunschweig.de/en/eis
--
-- Use of this source code is governed by an MIT-style
-- license that can be found in the LICENSE file or at
-- https://opensource.org/licenses/MIT.


package func_pkg is

  -- RTC
  constant FUNC_RTC_CNT_W_C : natural := 10;  -- Width of RTC counter
  
end package func_pkg;
